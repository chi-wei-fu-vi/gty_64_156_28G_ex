
package drp_reg_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
//  `include "reg_item_subscriber.svh"
  `include "vio_reg_block.svh"
  `include "gtye_channel_reg_block.svh"
  `include "gtye_common_reg_block.svh"
  `include "drp_top_reg_block.svh"
  `include "drp_reg_block.svh"
endpackage : drp_reg_pkg

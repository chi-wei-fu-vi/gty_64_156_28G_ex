package toplevel_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  import common_pkg::*;
  import common_env_pkg::*;
  import mm_pkg::*;
  typedef class toplevel_env;
  typedef class toplevel_config;
  `include "toplevel_env.svh"
  `include "toplevel_config.svh"
endpackage : toplevel_pkg
package toplevel_test_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  import common_pkg::*;
  import common_env_pkg::*;
  import toplevel_pkg::*;
  import mm_pkg::*;
  import drp_reg_pkg::*;
  typedef class base_test;
  typedef class seq_mm_item;
  `include "seq_examples.svh"
  `include "base_test.svh"
endpackage : toplevel_test_pkg
